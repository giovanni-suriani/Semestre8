library verilog;
use verilog.vl_types.all;
entity ReceptorTestbench is
end ReceptorTestbench;
