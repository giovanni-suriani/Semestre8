module PortaAND(entrada1,entrada2,saida);
input entrada1,entrada2;
output saida;
assign saida = entrada1 & entrada2;

endmodule

