library verilog;
use verilog.vl_types.all;
entity ProcessadorNrisc is
    port(
        clk             : in     vl_logic
    );
end ProcessadorNrisc;
