module somador(entrada1,entrada2,saida);
input[7:0] entrada1,entrada2;
output[7:0]  saida;

assign saida=entrada1+entrada2;


endmodule
