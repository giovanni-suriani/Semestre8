library verilog;
use verilog.vl_types.all;
entity SnoppingTestbench is
end SnoppingTestbench;
