library verilog;
use verilog.vl_types.all;
entity Memoryteste is
end Memoryteste;
